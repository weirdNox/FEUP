2018/19 - 2

.subckt ideal_op NonInv Inv Output Gain=100k
eE1 Output 0 NonInv Inv {Gain}
.ends

.subckt ideal_switch L R Phi
rS L R R=table(V(Phi), 0.5, 1000Meg, 0.8, 1)
.ends

vPhi1 Phi1 0 DC 0 PULSE(0 3 0                   2n 2n {DutyCycle*SamplingPeriod} {SamplingPeriod})
vPhi2 Phi2 0 DC 0 PULSE(0 3 {SamplingPeriod/2}  2n 2n {DutyCycle*SamplingPeriod} {SamplingPeriod})

.param C1 = 6p
.param C2 = 6p
.param Ca = 2p

.param SamplingFreq=50k
.param SamplingPeriod={1/SamplingFreq}
.param DutyCycle=.4

xS1    In     1      Phi1   ideal_switch
c1     1      2      {C1}
xS2    0      2      Phi1   ideal_switch
xS3    1      3      Phi2   ideal_switch
xS4    2      5      Phi2   ideal_switch
c2     5      0      {C2}
xS5    5      Out    Phi1   ideal_switch
xO     0      3      Out    ideal_op
cA     3      Out    {Ca}

xSB Out  OutS Phi1 ideal_switch
rO  OutS 0    5Meg

.param SignalFreq=3k
.param SignalPeriod={1/SignalFreq}
vIn In  0   SINE(0 1.5 {SignalFreq})
*vIn In  0   PULSE(0 1 {SignalPeriod/2} 1n 1n {SignalPeriod/2} {SignalPeriod})
.tran {3*SignalPeriod}
