* Switched Capacitor Filter

.subckt ideal_op NonInv Inv V+ V- Output Gain=100k
eE1 Output 0 NonInv Inv {Gain}
.ends

.subckt ideal_switch L R Phi
rS L R R=table(V(Phi), 0.5, 1000Meg, 0.8, 1)
.ends

vPhi1 Phi1 0 DC 0 PULSE(0 3 0                   2n 2n {DutyCycle*SamplingPeriod} {SamplingPeriod})
vPhi2 Phi2 0 DC 0 PULSE(0 3 {SamplingPeriod/2}  2n 2n {DutyCycle*SamplingPeriod} {SamplingPeriod})

* EXAMPLE
.param SamplingFreq=1Meg
.param SamplingPeriod={1/SamplingFreq}
.param DutyCycle=.4

xS1 In   2    Phi1 ideal_switch
xS2 2    0    Phi2 ideal_switch
c1  2    3    10p
xS3 3    0    Phi1 ideal_switch
xS4 3    4    Phi2 ideal_switch
c2  4    5    1p
xS5 5    Err  Phi1 ideal_switch
xS6 4    6    Phi1 ideal_switch
xS7 6    0    Phi2 ideal_switch
c3  6    7    0.5p
xS8 7    0    Phi2 ideal_switch
xS9 7    Out  Phi1 ideal_switch
xSA Out  5    Phi2 ideal_switch
xOp 0    4    0   0   Out ideal_op

xSB Out  OutS Phi1 ideal_switch
rO  OutS 0    5Meg

vE  Err  0    10

.param SignalFreq=25k
.param SignalPeriod={1/SignalFreq}
vIn In  0   SINE(0 1 {SignalFreq})
.tran {3*SignalPeriod}
